library ieee;
library work;
use work.components.all;
use ieee.std_logic_1164.all;

entity me_wb is
end entity;

architecture behavior of me_wb is
end architecture;
