library ieee;
library work;
use work.components.all;
use ieee.std_logic_1164.all;

entity ex_me is
end entity;

architecture behavior of ex_me is
end architecture;
