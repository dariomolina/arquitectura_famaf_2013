library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity problema_3_tb is
  generic (width : positive := 32);
end entity;

architecture test_bench of problema_3_tb is
  begin
end architecture;
