library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity problema_4_tb is
  generic (width : positive := 32);
end entity;

architecture test_bench of problema_4_tb is
  begin
end architecture;
