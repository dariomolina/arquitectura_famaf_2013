library ieee;
library work;
use ieee.std_logic_1164.all;
use work.components.all;

entity pipeline is
end entity;

architecture behavior of pipeline is
begin
end architecture;
